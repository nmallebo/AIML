    Mac OS X            	   2  �                                           ATTR        ,  �                 ,     com.apple.lastuseddate#PS      <   H  com.apple.macl     �  `  %com.apple.metadata:kMDItemWhereFroms   �     com.apple.provenance   �     com.apple.quarantine +�Hh    ��,     �Ma�L�����g ���P�Oܳ&��xՉ S����;MN�l��JL�                  bplist00�_https://files09.oaiusercontent.com/file-UnpreWNp97Ux1NwmHrREKW?se=2025-06-10T20%3A47%3A58Z&sp=r&sv=2024-08-04&sr=b&rscc=max-age%3D299%2C%20immutable%2C%20private&rscd=attachment%3B%20filename%3Disodata_cluster_multi_iter.sv&sig=9JP8XSS2Zh%2Biin4tr1IaJ6GvEhBA6wTbhvUW/7J5T9M%3D_https://chatgpt.com/  #                           : �3.i�-��q/0081;684898d2;Chrome; 