#######################################################################
####                                                               ####
####  The data contained in the file is created for educational    #### 
####  and training purposes only and are not recommended           ####
####  for fabrication                                              ####
####                                                               ####
#######################################################################
####                                                               ####
####  Copyright (C) 2013 Synopsys, Inc.                            ####
####                                                               ####
#######################################################################
####                                                               ####
####  The 32/28nm Generic Library ("Library") is unsupported       ####    
####  Confidential Information of Synopsys, Inc. ("Synopsys")      ####    
####  provided to you as Documentation under the terms of the      ####    
####  End User Software License Agreement between you or your      ####    
####  employer and Synopsys ("License Agreement") and you agree    ####    
####  not to distribute or disclose the Library without the        ####    
####  prior written consent of Synopsys. The Library IS NOT an     ####    
####  item of Licensed Software or Licensed Product under the      ####    
####  License Agreement.  Synopsys and/or its licensors own        ####    
####  and shall retain all right, title and interest in and        ####    
####  to the Library and all modifications thereto, including      ####    
####  all intellectual property rights embodied therein. All       ####    
####  rights in and to any Library modifications you make are      ####    
####  hereby assigned to Synopsys. If you do not agree with        ####    
####  this notice, including the disclaimer below, then you        ####    
####  are not authorized to use the Library.                       ####    
####                                                               ####  
####                                                               ####      
####  THIS LIBRARY IS BEING DISTRIBUTED BY SYNOPSYS SOLELY ON AN   ####
####  "AS IS" BASIS, WITH NO INTELLECUTAL PROPERTY                 ####
####  INDEMNIFICATION AND NO SUPPORT. ANY EXPRESS OR IMPLIED       ####
####  WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED       ####
####  WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR   ####
####  PURPOSE ARE HEREBY DISCLAIMED. IN NO EVENT SHALL SYNOPSYS    ####
####  BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     ####
####  EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT      ####
####  LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;     ####
####  LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)     ####
####  HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN    ####
####  CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE    ####
####  OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS      ####
####  DOCUMENTATION, EVEN IF ADVISED OF THE POSSIBILITY OF         ####
####  SUCH DAMAGE.                                                 #### 
####                                                               ####  
#######################################################################

# 
# LEF OUT 
# User Name : edbab 
# Date : Mon Dec 24 17:39:17 2012
# 
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;

MACRO PLL
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 113.223 BY 48.108 ;
  SYMMETRY X Y R90 ;

  PIN AVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 94.6080 47.7650 95.1080 48.1080 ;
    END
    ANTENNADIFFAREA 42.2555 LAYER M6 ;
    ANTENNADIFFAREA 42.2555 LAYER M7 ;
    ANTENNADIFFAREA 42.2555 LAYER M8 ;
    ANTENNADIFFAREA 42.2555 LAYER M9 ;
    ANTENNADIFFAREA 42.2555 LAYER MRDL ;
    ANTENNAGATEAREA 0.322 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 19.7555 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 19.7555 LAYER M6 ;
    ANTENNAMAXAREACAR 94.42332 LAYER M6 ;
    ANTENNAGATEAREA 0.322 LAYER M7 ;
    ANTENNAGATEAREA 0.322 LAYER M8 ;
    ANTENNAGATEAREA 0.322 LAYER M9 ;
    ANTENNAGATEAREA 0.322 LAYER MRDL ;
  END AVDD

  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M6 ;
        RECT 101.9890 47.8690 102.4890 48.1080 ;
    END
    ANTENNADIFFAREA 19.75664 LAYER M6 ;
    ANTENNADIFFAREA 19.75664 LAYER M7 ;
    ANTENNADIFFAREA 19.75664 LAYER M8 ;
    ANTENNADIFFAREA 19.75664 LAYER M9 ;
    ANTENNADIFFAREA 19.75664 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 21.4715 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 21.4715 LAYER M6 ;
  END DVDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M6 ;
        RECT 107.3470 47.8800 107.8470 48.1080 ;
    END
    ANTENNADIFFAREA 285.3474 LAYER M6 ;
    ANTENNADIFFAREA 285.3474 LAYER M7 ;
    ANTENNADIFFAREA 285.3474 LAYER M8 ;
    ANTENNADIFFAREA 285.3474 LAYER M9 ;
    ANTENNADIFFAREA 285.3474 LAYER MRDL ;
    ANTENNAGATEAREA 0.84 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 22.283 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 22.283 LAYER M6 ;
    ANTENNAMAXAREACAR 78.7198 LAYER M6 ;
    ANTENNAGATEAREA 0.84 LAYER M7 ;
    ANTENNAGATEAREA 0.84 LAYER M8 ;
    ANTENNAGATEAREA 0.84 LAYER M9 ;
    ANTENNAGATEAREA 0.84 LAYER MRDL ;
  END VSS

  PIN PLL_BYPASS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.0950 29.0860 113.2230 29.2770 ;
    END
    ANTENNAGATEAREA 0.144 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
    ANTENNAMAXAREACAR 17.46132 LAYER M6 ;
    ANTENNAGATEAREA 0.144 LAYER M7 ;
    ANTENNAGATEAREA 0.144 LAYER M8 ;
    ANTENNAGATEAREA 0.144 LAYER M9 ;
    ANTENNAGATEAREA 0.144 LAYER MRDL ;
  END PLL_BYPASS

  PIN CLK_1X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.0860 23.4830 113.2230 23.6740 ;
    END
    ANTENNADIFFAREA 0.12934 LAYER M6 ;
    ANTENNADIFFAREA 0.12934 LAYER M7 ;
    ANTENNADIFFAREA 0.12934 LAYER M8 ;
    ANTENNADIFFAREA 0.12934 LAYER M9 ;
    ANTENNADIFFAREA 0.12934 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
  END CLK_1X

  PIN CLK_2X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.0860 21.7560 113.2230 21.9470 ;
    END
    ANTENNADIFFAREA 0.12934 LAYER M6 ;
    ANTENNADIFFAREA 0.12934 LAYER M7 ;
    ANTENNADIFFAREA 0.12934 LAYER M8 ;
    ANTENNADIFFAREA 0.12934 LAYER M9 ;
    ANTENNADIFFAREA 0.12934 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
  END CLK_2X

  PIN REF_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.0880 12.6490 113.2230 12.8400 ;
    END
    ANTENNAGATEAREA 0.096 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
    ANTENNAMAXAREACAR 29.39242 LAYER M6 ;
    ANTENNAGATEAREA 0.096 LAYER M7 ;
    ANTENNAGATEAREA 0.096 LAYER M8 ;
    ANTENNAGATEAREA 0.096 LAYER M9 ;
    ANTENNAGATEAREA 0.096 LAYER MRDL ;
  END REF_CLK

  PIN FB_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 87.2850 0.0000 87.4760 0.1260 ;
    END
    ANTENNAGATEAREA 0.024 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
    ANTENNAMAXAREACAR 27.84097 LAYER M6 ;
    ANTENNAGATEAREA 0.024 LAYER M7 ;
    ANTENNAGATEAREA 0.024 LAYER M8 ;
    ANTENNAGATEAREA 0.024 LAYER M9 ;
    ANTENNAGATEAREA 0.024 LAYER MRDL ;
  END FB_CLK

  PIN FB_MODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 88.5390 0.0000 88.7300 0.1270 ;
    END
    ANTENNAGATEAREA 0.048 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
    ANTENNAMAXAREACAR 12.95897 LAYER M6 ;
    ANTENNAGATEAREA 0.048 LAYER M7 ;
    ANTENNAGATEAREA 0.048 LAYER M8 ;
    ANTENNAGATEAREA 0.048 LAYER M9 ;
    ANTENNAGATEAREA 0.048 LAYER MRDL ;
  END FB_MODE

  PIN CLK_4X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 113.0800 20.0160 113.2230 20.2070 ;
    END
    ANTENNADIFFAREA 0.12934 LAYER M6 ;
    ANTENNADIFFAREA 0.12934 LAYER M7 ;
    ANTENNADIFFAREA 0.12934 LAYER M8 ;
    ANTENNADIFFAREA 0.12934 LAYER M9 ;
    ANTENNADIFFAREA 0.12934 LAYER MRDL ;
    ANTENNAPARTIALMETALAREA 0.081366 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 0.081366 LAYER M6 ;
  END CLK_4X
  OBS
    LAYER MRDL ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M6 ;
      RECT 87.5320 29.3330 88.4830 47.7090 ;
      RECT 0.0000 29.3330 87.2290 47.7090 ;
      RECT 112.7970 29.0300 113.0240 29.0860 ;
      RECT 112.7970 12.5930 113.0240 12.8960 ;
      RECT 112.7970 29.2770 113.0240 29.3330 ;
      RECT 112.7970 29.0860 113.0310 29.2770 ;
      RECT 87.5320 0.1900 88.4750 0.1910 ;
      RECT 87.5400 0.1830 88.4750 0.1900 ;
      RECT 94.6080 12.5930 95.1080 12.8960 ;
      RECT 94.6080 29.0300 95.1080 29.3330 ;
      RECT 101.9890 12.5930 102.4890 12.8960 ;
      RECT 101.9890 47.7090 102.4890 47.7590 ;
      RECT 101.9890 29.0300 102.4890 29.3330 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 12.5930 107.8470 12.8960 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 29.0300 107.8470 29.3330 ;
      RECT 107.3470 47.7090 107.8470 47.7700 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 107.3470 21.7000 107.8470 23.7380 ;
      RECT 94.6080 21.7000 95.1080 23.4270 ;
      RECT 94.6080 23.4190 95.1080 23.7300 ;
      RECT 94.6080 19.9600 95.1080 20.2710 ;
      RECT 94.6080 23.4190 95.1080 23.7300 ;
      RECT 94.6080 19.9600 95.1080 20.2710 ;
      RECT 94.6080 21.7000 95.1080 23.4270 ;
      RECT 101.9890 21.7000 102.4890 23.4270 ;
      RECT 101.9890 19.9600 102.4890 20.2710 ;
      RECT 101.9890 23.4190 102.4890 23.7300 ;
      RECT 101.9890 23.4190 102.4890 23.7300 ;
      RECT 101.9890 19.9600 102.4890 20.2710 ;
      RECT 101.9890 21.7000 102.4890 23.4270 ;
      RECT 112.7970 21.7000 113.0220 23.4270 ;
      RECT 112.7970 21.7000 113.0220 23.7300 ;
      RECT 112.7970 21.7000 113.0220 23.4270 ;
      RECT 112.7970 21.7000 113.0220 23.7300 ;
      RECT 87.2290 0.1900 88.4750 0.1910 ;
      RECT 87.2290 0.1910 91.7870 0.4260 ;
      RECT 87.5320 0.4260 88.4830 12.5930 ;
      RECT 88.7860 23.4190 113.0220 23.4270 ;
      RECT 88.7860 21.6920 113.0220 21.7000 ;
      RECT 88.7860 20.2630 113.0160 20.2710 ;
      RECT 88.7860 0.4260 91.7870 8.5970 ;
      RECT 88.7860 22.0030 113.0220 22.0110 ;
      RECT 88.7860 20.2710 113.0240 21.6920 ;
      RECT 88.7860 22.0110 113.0240 23.4190 ;
      RECT 88.7860 16.9590 113.0160 19.9600 ;
      RECT 88.7860 23.7300 113.0220 26.7310 ;
      RECT 101.9890 47.4580 102.4890 47.7590 ;
      RECT 107.3470 19.9600 107.8470 20.2630 ;
      RECT 112.7970 19.9600 113.0160 20.2630 ;
      RECT 112.7970 29.0300 113.0240 29.3330 ;
      RECT 88.7860 29.3330 94.4980 47.7090 ;
      RECT 88.7860 29.3330 94.4980 47.7090 ;
      RECT 88.7860 47.6550 94.4980 47.7090 ;
      RECT 95.1640 0.1830 101.9330 8.5970 ;
      RECT 95.1640 0.1830 101.9330 5.1650 ;
      RECT 88.7860 29.3330 113.0240 47.6550 ;
      RECT 95.2180 47.6550 113.0240 47.7090 ;
      RECT 95.2180 29.3330 113.0240 47.7090 ;
      RECT 95.2180 29.3330 113.0240 47.7090 ;
      RECT 102.5450 0.1830 107.2910 8.5970 ;
      RECT 102.5450 0.1830 107.2910 3.5420 ;
      RECT 95.1640 5.1650 113.0240 8.5970 ;
      RECT 102.5450 3.5420 113.0240 8.5970 ;
      RECT 102.5450 3.5420 113.0240 5.1650 ;
      RECT 107.9030 0.1830 113.0240 8.5970 ;
      RECT 107.9030 0.1830 113.0240 3.5420 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1830 87.2210 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1830 87.2210 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1830 87.2210 12.5930 ;
      RECT 0.0000 0.1830 87.2210 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 0.0000 0.1830 87.2210 12.5930 ;
      RECT 0.0000 0.1900 87.2290 12.5930 ;
      RECT 88.7860 8.5970 113.0240 12.5930 ;
      RECT 88.7940 0.1830 94.5520 8.5970 ;
      RECT 88.7940 0.1830 94.5520 8.5970 ;
      RECT 88.7940 0.1830 94.5520 8.5970 ;
      RECT 88.7860 23.7380 113.0240 29.0300 ;
      RECT 88.7860 12.8960 113.0240 19.9520 ;
      RECT 87.5320 23.7300 88.4830 29.0300 ;
      RECT 0.0000 23.7300 87.2290 29.0300 ;
      RECT 87.5320 22.0030 88.4830 23.4270 ;
      RECT 0.0000 22.0030 87.2290 23.4270 ;
      RECT 87.5320 20.2630 88.4830 21.7000 ;
      RECT 0.0000 20.2630 87.2290 21.7000 ;
      RECT 87.5320 12.8960 88.4830 19.9600 ;
      RECT 0.0000 12.8960 87.2290 19.9600 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M3 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER M1 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER PO ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
    LAYER CO ;
      RECT 0.0000 0.0000 113.2230 48.1080 ;
  END
END PLL
  
END LIBRARY
