    Mac OS X            	   2  �     �                                      ATTR      �    �                    H  com.apple.macl     L  g  %com.apple.metadata:kMDItemWhereFroms   �     com.apple.provenance   �     com.apple.quarantine  �Ma�L�����g ���P�Oܳ&��xՉ S����;MN�l��JL�                  bplist00�_https://files.oaiusercontent.com/file-Prw6HneHvRPVtJN5G5B1wa?se=2025-06-10T22%3A40%3A32Z&sp=r&sv=2024-08-04&sr=b&rscc=max-age%3D299%2C%20immutable%2C%20private&rscd=attachment%3B%20filename%3Dtb_isodata_cluster_scaled_real_output.sv&sig=El5KfOzI1mbE3epQ8cfO0ry9OQwBQUFFF7tvKnPMygI%3D_https://chatgpt.com/  *                           A �3.i�-��q/0081;6848b334;Chrome; 